`ifndef COLOR_SVH
`define COLOR_SVH

`define BLACK_COLOR $write("\033[30m");
`define RED_COLOR $write("\033[31m");
`define GREEN_COLOR $write("\033[32m");
`define YELLOW_COLOR $write("\033[33m");
`define BLUE_COLOR $write("\033[34m");
`define MAGENTA_COLOR $write("\033[35m");
`define CYAN_COLOR $write("\033[36m");
`define WHITE_COLOR $write("\033[37m");
`define GRAY_COLOR $write("\033[90m");
`define RESET_COLOR $write("\033[0m");

`endif
